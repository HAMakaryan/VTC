module ch4_test;



endmodule
