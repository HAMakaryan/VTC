//    file 06_05_03_Ripple_Counter.v

module 06_05_03_Ripple_Counter(

);


endmodule
