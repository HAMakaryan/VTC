module ripple_adder_top;

//Draft


#(
// Parameter Declaration. This can be redefined
  .N = 16 // 4-bit bus by default
)
uq
(
  .co   (lalsjalksj),
  .sum  (lalsjalksj),
  .a0   (lalsjalksj),
  .a1   (lalsjalksj),
  .ci
);



#(
// Parameter Declaration. This can be redefined
  .N = 32 // 4-bit bus by default
)
u2
(
  .co   (lalsjalksj),
  .sum  (lalsjalksj),
  .a0   (lalsjalksj),
  .a1   (lalsjalksj),
  .ci
);





endmodule
