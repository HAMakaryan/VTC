module lcd_top;



endmodule

